/* arachne-pnr 0.1+20180513git5d830dd (git sha1 5d830dd, g++ 9.3.0-6ubuntu1 -O2 -fdebug-prefix-map=/build/arachne-pnr-AaC6iz/arachne-pnr-0.1+20180513git5d830dd=. -fstack-protector-strong -O2 -DNDEBUG) */
module top(input CLK, output VGA_HS, output VGA_VS, output VGA_R0, output VGA_R1, output VGA_R2, output VGA_G0, output VGA_G1, output VGA_G2, output VGA_B0, output VGA_B1, output VGA_B2);
  wire \$abc$1026$auto$alumacc.cc:474:replace_alu$92.BB[0] ;
  wire \$abc$1026$auto$alumacc.cc:474:replace_alu$92.BB[1] ;
  wire \$abc$1026$auto$alumacc.cc:474:replace_alu$92.BB[2] ;
  wire \$abc$1026$auto$alumacc.cc:474:replace_alu$92.BB[3] ;
  wire \$abc$1026$auto$alumacc.cc:474:replace_alu$92.BB[4] ;
  wire \$abc$1026$auto$alumacc.cc:474:replace_alu$92.BB[5] ;
  wire \$abc$1026$auto$alumacc.cc:474:replace_alu$92.BB[6] ;
  wire \$abc$1026$auto$alumacc.cc:474:replace_alu$92.BB[7] ;
  wire \$abc$1026$auto$alumacc.cc:474:replace_alu$92.BB[8] ;
  wire \$abc$1026$auto$dff2dffe.cc:175:make_patterns_logic$868 ;
  wire \$abc$1026$auto$simplemap.cc:127:simplemap_reduce$263[0]_new_inv_ ;
  wire \$abc$1026$auto$simplemap.cc:127:simplemap_reduce$310[0]_new_inv_ ;
  wire $abc$1026$new_n100_;
  wire $abc$1026$new_n103_;
  wire $abc$1026$new_n108_;
  wire $abc$1026$new_n109_;
  wire $abc$1026$new_n110_;
  wire $abc$1026$new_n117_;
  wire $abc$1026$new_n118_;
  wire $abc$1026$new_n69_;
  wire $abc$1026$new_n72_;
  wire $abc$1026$new_n73_;
  wire $abc$1026$new_n97_;
  wire $abc$1026$new_n98_;
  wire $abc$1026$new_n99_;
  wire $abc$1026$visible_new_;
  wire \$auto$alumacc.cc:474:replace_alu$104.C[2] ;
  wire \$auto$alumacc.cc:474:replace_alu$104.C[3] ;
  wire \$auto$alumacc.cc:474:replace_alu$104.C[4] ;
  wire \$auto$alumacc.cc:474:replace_alu$104.C[5] ;
  wire \$auto$alumacc.cc:474:replace_alu$104.C[6] ;
  wire \$auto$alumacc.cc:474:replace_alu$104.C[7] ;
  wire \$auto$alumacc.cc:474:replace_alu$104.C[8] ;
  wire \$auto$alumacc.cc:474:replace_alu$104.C[9] ;
  wire \$auto$alumacc.cc:474:replace_alu$92.C[1] ;
  wire \$auto$alumacc.cc:474:replace_alu$92.C[2] ;
  wire \$auto$alumacc.cc:474:replace_alu$92.C[3] ;
  wire \$auto$alumacc.cc:474:replace_alu$92.C[4] ;
  wire \$auto$alumacc.cc:474:replace_alu$92.C[5] ;
  wire \$auto$alumacc.cc:474:replace_alu$92.C[6] ;
  wire \$auto$alumacc.cc:474:replace_alu$92.C[7] ;
  wire \$auto$alumacc.cc:474:replace_alu$92.C[8] ;
  wire \$auto$alumacc.cc:474:replace_alu$95.C[10] ;
  wire \$auto$alumacc.cc:474:replace_alu$95.C[11] ;
  wire \$auto$alumacc.cc:474:replace_alu$95.C[12] ;
  wire \$auto$alumacc.cc:474:replace_alu$95.C[13] ;
  wire \$auto$alumacc.cc:474:replace_alu$95.C[14] ;
  wire \$auto$alumacc.cc:474:replace_alu$95.C[15] ;
  wire \$auto$alumacc.cc:474:replace_alu$95.C[16] ;
  wire \$auto$alumacc.cc:474:replace_alu$95.C[17] ;
  wire \$auto$alumacc.cc:474:replace_alu$95.C[18] ;
  wire \$auto$alumacc.cc:474:replace_alu$95.C[19] ;
  wire \$auto$alumacc.cc:474:replace_alu$95.C[20] ;
  wire \$auto$alumacc.cc:474:replace_alu$95.C[21] ;
  wire \$auto$alumacc.cc:474:replace_alu$95.C[22] ;
  wire \$auto$alumacc.cc:474:replace_alu$95.C[23] ;
  wire \$auto$alumacc.cc:474:replace_alu$95.C[24] ;
  wire \$auto$alumacc.cc:474:replace_alu$95.C[25] ;
  wire \$auto$alumacc.cc:474:replace_alu$95.C[26] ;
  wire \$auto$alumacc.cc:474:replace_alu$95.C[27] ;
  wire \$auto$alumacc.cc:474:replace_alu$95.C[28] ;
  wire \$auto$alumacc.cc:474:replace_alu$95.C[2] ;
  wire \$auto$alumacc.cc:474:replace_alu$95.C[3] ;
  wire \$auto$alumacc.cc:474:replace_alu$95.C[4] ;
  wire \$auto$alumacc.cc:474:replace_alu$95.C[5] ;
  wire \$auto$alumacc.cc:474:replace_alu$95.C[6] ;
  wire \$auto$alumacc.cc:474:replace_alu$95.C[7] ;
  wire \$auto$alumacc.cc:474:replace_alu$95.C[8] ;
  wire \$auto$alumacc.cc:474:replace_alu$95.C[9] ;
  wire \$auto$alumacc.cc:474:replace_alu$98.C[2] ;
  wire \$auto$alumacc.cc:474:replace_alu$98.C[3] ;
  wire \$auto$alumacc.cc:474:replace_alu$98.C[4] ;
  wire \$auto$alumacc.cc:474:replace_alu$98.C[5] ;
  wire \$auto$alumacc.cc:474:replace_alu$98.C[6] ;
  wire \$auto$alumacc.cc:474:replace_alu$98.C[7] ;
  wire \$auto$alumacc.cc:474:replace_alu$98.C[8] ;
  wire \$auto$alumacc.cc:474:replace_alu$98.C[9] ;
  wire $false = 0;
  wire $true = 1;
  wire CLK$2;
  wire VGA_B0$2;
  wire VGA_B1$2;
  wire VGA_B2$2;
  wire VGA_G0$2;
  wire VGA_G1$2;
  wire VGA_G2$2;
  wire VGA_HS$2;
  wire VGA_R0$2;
  wire VGA_R1$2;
  wire VGA_R2$2;
  wire VGA_VS$2;
  wire \in_b[0] ;
  wire \in_b[1] ;
  wire \in_b[2] ;
  wire \in_g[0] ;
  wire \in_g[1] ;
  wire \in_g[2] ;
  wire \in_r[0] ;
  wire \in_r[1] ;
  wire \in_r[2] ;
  wire \ra_time[0] ;
  wire \ra_time[0]$2 ;
  wire \ra_time[10] ;
  wire \ra_time[11] ;
  wire \ra_time[12] ;
  wire \ra_time[13] ;
  wire \ra_time[14] ;
  wire \ra_time[15] ;
  wire \ra_time[16] ;
  wire \ra_time[17] ;
  wire \ra_time[18] ;
  wire \ra_time[19] ;
  wire \ra_time[1] ;
  wire \ra_time[20] ;
  wire \ra_time[21] ;
  wire \ra_time[22] ;
  wire \ra_time[23] ;
  wire \ra_time[24] ;
  wire \ra_time[25] ;
  wire \ra_time[26] ;
  wire \ra_time[27] ;
  wire \ra_time[28] ;
  wire \ra_time[2] ;
  wire \ra_time[3] ;
  wire \ra_time[4] ;
  wire \ra_time[5] ;
  wire \ra_time[6] ;
  wire \ra_time[7] ;
  wire \ra_time[8] ;
  wire \ra_time[9] ;
  wire \uut.vga_h_pixel_tracker.o_reset_counter ;
  wire \uut.vga_h_pixel_tracker.ra_coord[0] ;
  wire \uut.vga_h_pixel_tracker.ra_coord[0]$2 ;
  wire \uut.vga_h_pixel_tracker.ra_coord[1] ;
  wire \uut.vga_h_pixel_tracker.ra_coord[2] ;
  wire \uut.vga_h_pixel_tracker.ra_coord[3] ;
  wire \uut.vga_h_pixel_tracker.ra_coord[4] ;
  wire \uut.vga_h_pixel_tracker.ra_coord[5] ;
  wire \uut.vga_h_pixel_tracker.ra_coord[6] ;
  wire \uut.vga_h_pixel_tracker.ra_coord[7] ;
  wire \uut.vga_h_pixel_tracker.ra_coord[8] ;
  wire \uut.vga_h_pixel_tracker.ra_coord[9] ;
  wire \uut.vga_h_pixel_tracker.ra_state[0] ;
  wire \uut.vga_h_pixel_tracker.ra_state[1] ;
  wire \uut.vga_v_pixel_tracker.o_reset_counter ;
  wire \uut.vga_v_pixel_tracker.ra_coord[0] ;
  wire \uut.vga_v_pixel_tracker.ra_coord[0]$2 ;
  wire \uut.vga_v_pixel_tracker.ra_coord[1] ;
  wire \uut.vga_v_pixel_tracker.ra_coord[2] ;
  wire \uut.vga_v_pixel_tracker.ra_coord[3] ;
  wire \uut.vga_v_pixel_tracker.ra_coord[4] ;
  wire \uut.vga_v_pixel_tracker.ra_coord[5] ;
  wire \uut.vga_v_pixel_tracker.ra_coord[6] ;
  wire \uut.vga_v_pixel_tracker.ra_coord[7] ;
  wire \uut.vga_v_pixel_tracker.ra_coord[8] ;
  wire \uut.vga_v_pixel_tracker.ra_coord[9] ;
  wire \uut.vga_v_pixel_tracker.ra_state[0] ;
  wire \uut.vga_v_pixel_tracker.ra_state[1] ;
  SB_IO #(
    .PIN_TYPE(6'b000001)
  ) $inst0 (
    .PACKAGE_PIN(CLK),
    .D_IN_0(CLK$2)
  );
  SB_IO #(
    .PIN_TYPE(6'b011001)
  ) $inst1 (
    .PACKAGE_PIN(VGA_B0),
    .D_OUT_0(VGA_B0$2)
  );
  SB_IO #(
    .PIN_TYPE(6'b011001)
  ) $inst2 (
    .PACKAGE_PIN(VGA_B1),
    .D_OUT_0(VGA_B1$2)
  );
  SB_IO #(
    .PIN_TYPE(6'b011001)
  ) $inst3 (
    .PACKAGE_PIN(VGA_B2),
    .D_OUT_0(VGA_B2$2)
  );
  SB_IO #(
    .PIN_TYPE(6'b011001)
  ) $inst4 (
    .PACKAGE_PIN(VGA_G0),
    .D_OUT_0(VGA_G0$2)
  );
  SB_IO #(
    .PIN_TYPE(6'b011001)
  ) $inst5 (
    .PACKAGE_PIN(VGA_G1),
    .D_OUT_0(VGA_G1$2)
  );
  SB_IO #(
    .PIN_TYPE(6'b011001)
  ) $inst6 (
    .PACKAGE_PIN(VGA_G2),
    .D_OUT_0(VGA_G2$2)
  );
  SB_IO #(
    .PIN_TYPE(6'b011001)
  ) $inst7 (
    .PACKAGE_PIN(VGA_HS),
    .D_OUT_0(VGA_HS$2)
  );
  SB_IO #(
    .PIN_TYPE(6'b011001)
  ) $inst8 (
    .PACKAGE_PIN(VGA_R0),
    .D_OUT_0(VGA_R0$2)
  );
  SB_IO #(
    .PIN_TYPE(6'b011001)
  ) $inst9 (
    .PACKAGE_PIN(VGA_R1),
    .D_OUT_0(VGA_R1$2)
  );
  SB_IO #(
    .PIN_TYPE(6'b011001)
  ) $inst10 (
    .PACKAGE_PIN(VGA_R2),
    .D_OUT_0(VGA_R2$2)
  );
  SB_IO #(
    .PIN_TYPE(6'b011001)
  ) $inst11 (
    .PACKAGE_PIN(VGA_VS),
    .D_OUT_0(VGA_VS$2)
  );
  (* src="top.v:85|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:86|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0101101010100101)
  ) $inst12 (
    .I0($false),
    .I1($false),
    .I2(\ra_time[0] ),
    .I3($false),
    .CLK(CLK$2),
    .CEN($true),
    .SR($false),
    .O(\ra_time[0] )
  );
  (* src="top.v:85|/usr/bin/../share/yosys/ice40/cells_map.v:8|/usr/bin/../share/yosys/ice40/cells_map.v:40" *)
  ICESTORM_LC #(
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(2'b01)
  ) $inst13 (
    .I0(\ra_time[1] ),
    .I1($false),
    .I2($false),
    .I3($false),
    .CLK(CLK$2),
    .CEN(\ra_time[0] ),
    .SR($false),
    .O(\ra_time[1] )
  );
  (* src="top.v:85|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:86|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst14 (
    .I0($false),
    .I1($false),
    .I2(\ra_time[2] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$95.C[2] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$95.C[2] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR($false),
    .O(\ra_time[2] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$95.C[3] )
  );
  (* src="top.v:85|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:86|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst15 (
    .I0($false),
    .I1($false),
    .I2(\ra_time[3] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$95.C[3] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$95.C[3] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR($false),
    .O(\ra_time[3] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$95.C[4] )
  );
  (* src="top.v:85|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:86|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst16 (
    .I0($false),
    .I1($false),
    .I2(\ra_time[4] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$95.C[4] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$95.C[4] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR($false),
    .O(\ra_time[4] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$95.C[5] )
  );
  (* src="top.v:85|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:86|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst17 (
    .I0($false),
    .I1($false),
    .I2(\ra_time[5] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$95.C[5] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$95.C[5] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR($false),
    .O(\ra_time[5] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$95.C[6] )
  );
  (* src="top.v:85|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:86|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst18 (
    .I0($false),
    .I1($false),
    .I2(\ra_time[6] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$95.C[6] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$95.C[6] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR($false),
    .O(\ra_time[6] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$95.C[7] )
  );
  (* src="top.v:85|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:86|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst19 (
    .I0($false),
    .I1($false),
    .I2(\ra_time[7] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$95.C[7] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$95.C[7] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR($false),
    .O(\ra_time[7] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$95.C[8] )
  );
  (* src="top.v:85|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:86|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst20 (
    .I0($false),
    .I1($false),
    .I2(\ra_time[8] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$95.C[8] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$95.C[8] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR($false),
    .O(\ra_time[8] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$95.C[9] )
  );
  (* src="top.v:85|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:86|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst21 (
    .I0($false),
    .I1($false),
    .I2(\ra_time[9] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$95.C[9] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$95.C[9] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR($false),
    .O(\ra_time[9] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$95.C[10] )
  );
  (* src="top.v:85|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:86|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst22 (
    .I0($false),
    .I1($false),
    .I2(\ra_time[10] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$95.C[10] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$95.C[10] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR($false),
    .O(\ra_time[10] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$95.C[11] )
  );
  (* src="top.v:85|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:86|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst23 (
    .I0($false),
    .I1($false),
    .I2(\ra_time[11] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$95.C[11] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$95.C[11] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR($false),
    .O(\ra_time[11] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$95.C[12] )
  );
  (* src="top.v:85|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:86|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst24 (
    .I0($false),
    .I1($false),
    .I2(\ra_time[12] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$95.C[12] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$95.C[12] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR($false),
    .O(\ra_time[12] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$95.C[13] )
  );
  (* src="top.v:85|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:86|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst25 (
    .I0($false),
    .I1($false),
    .I2(\ra_time[13] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$95.C[13] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$95.C[13] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR($false),
    .O(\ra_time[13] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$95.C[14] )
  );
  (* src="top.v:85|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:86|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst26 (
    .I0($false),
    .I1($false),
    .I2(\ra_time[14] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$95.C[14] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$95.C[14] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR($false),
    .O(\ra_time[14] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$95.C[15] )
  );
  (* src="top.v:85|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:86|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst27 (
    .I0($false),
    .I1($false),
    .I2(\ra_time[15] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$95.C[15] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$95.C[15] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR($false),
    .O(\ra_time[15] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$95.C[16] )
  );
  (* src="top.v:85|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:86|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst28 (
    .I0($false),
    .I1($false),
    .I2(\ra_time[16] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$95.C[16] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$95.C[16] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR($false),
    .O(\ra_time[16] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$95.C[17] )
  );
  (* src="top.v:85|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:86|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst29 (
    .I0($false),
    .I1($false),
    .I2(\ra_time[17] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$95.C[17] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$95.C[17] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR($false),
    .O(\ra_time[17] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$95.C[18] )
  );
  (* src="top.v:85|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:86|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst30 (
    .I0($false),
    .I1($false),
    .I2(\ra_time[18] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$95.C[18] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$95.C[18] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR($false),
    .O(\ra_time[18] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$95.C[19] )
  );
  (* src="top.v:85|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:86|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst31 (
    .I0($false),
    .I1($false),
    .I2(\ra_time[19] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$95.C[19] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$95.C[19] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR($false),
    .O(\ra_time[19] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$95.C[20] )
  );
  (* src="top.v:85|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:86|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst32 (
    .I0($false),
    .I1($false),
    .I2(\ra_time[20] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$95.C[20] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$95.C[20] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR($false),
    .O(\ra_time[20] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$95.C[21] )
  );
  (* src="top.v:85|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:86|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst33 (
    .I0($false),
    .I1($false),
    .I2(\ra_time[21] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$95.C[21] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$95.C[21] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR($false),
    .O(\ra_time[21] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$95.C[22] )
  );
  (* src="top.v:85|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:86|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst34 (
    .I0($false),
    .I1($false),
    .I2(\ra_time[22] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$95.C[22] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$95.C[22] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR($false),
    .O(\ra_time[22] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$95.C[23] )
  );
  (* src="top.v:85|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:86|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst35 (
    .I0($false),
    .I1($false),
    .I2(\ra_time[23] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$95.C[23] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$95.C[23] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR($false),
    .O(\ra_time[23] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$95.C[24] )
  );
  (* src="top.v:85|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:86|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst36 (
    .I0($false),
    .I1($false),
    .I2(\ra_time[24] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$95.C[24] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$95.C[24] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR($false),
    .O(\ra_time[24] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$95.C[25] )
  );
  (* src="top.v:85|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:86|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst37 (
    .I0($false),
    .I1($false),
    .I2(\ra_time[25] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$95.C[25] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$95.C[25] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR($false),
    .O(\ra_time[25] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$95.C[26] )
  );
  (* src="top.v:85|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:86|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst38 (
    .I0($false),
    .I1($false),
    .I2(\ra_time[26] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$95.C[26] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$95.C[26] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR($false),
    .O(\ra_time[26] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$95.C[27] )
  );
  (* src="top.v:85|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:86|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst39 (
    .I0($false),
    .I1($false),
    .I2(\ra_time[27] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$95.C[27] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$95.C[27] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR($false),
    .O(\ra_time[27] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$95.C[28] )
  );
  (* src="top.v:85|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:86|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst40 (
    .I0($false),
    .I1($false),
    .I2(\ra_time[28] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$95.C[28] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR($false),
    .O(\ra_time[28] )
  );
  (* src="top.v:60|../../../lib/interface/Vga.v:88|../../../lib/interface/Vga.v:42|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:60|../../../lib/interface/Vga.v:88|../../../lib/interface/Vga.v:44|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0101101010100101)
  ) $inst41 (
    .I0($false),
    .I1($false),
    .I2(\uut.vga_h_pixel_tracker.ra_coord[0] ),
    .I3($false),
    .CLK(CLK$2),
    .CEN($true),
    .SR(\uut.vga_h_pixel_tracker.o_reset_counter ),
    .O(\uut.vga_h_pixel_tracker.ra_coord[0] )
  );
  (* src="top.v:60|../../../lib/interface/Vga.v:88|../../../lib/interface/Vga.v:42|/usr/bin/../share/yosys/ice40/cells_map.v:8|/usr/bin/../share/yosys/ice40/cells_map.v:40" *)
  ICESTORM_LC #(
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(2'b01)
  ) $inst42 (
    .I0(\uut.vga_h_pixel_tracker.ra_coord[1] ),
    .I1($false),
    .I2($false),
    .I3($false),
    .CLK(CLK$2),
    .CEN(\uut.vga_h_pixel_tracker.ra_coord[0] ),
    .SR(\uut.vga_h_pixel_tracker.o_reset_counter ),
    .O(\uut.vga_h_pixel_tracker.ra_coord[1] )
  );
  (* src="top.v:60|../../../lib/interface/Vga.v:88|../../../lib/interface/Vga.v:42|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:60|../../../lib/interface/Vga.v:88|../../../lib/interface/Vga.v:44|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst43 (
    .I0($false),
    .I1($false),
    .I2(\uut.vga_h_pixel_tracker.ra_coord[2] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$98.C[2] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$98.C[2] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR(\uut.vga_h_pixel_tracker.o_reset_counter ),
    .O(\uut.vga_h_pixel_tracker.ra_coord[2] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$98.C[3] )
  );
  (* src="top.v:60|../../../lib/interface/Vga.v:88|../../../lib/interface/Vga.v:42|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:60|../../../lib/interface/Vga.v:88|../../../lib/interface/Vga.v:44|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst44 (
    .I0($false),
    .I1($false),
    .I2(\uut.vga_h_pixel_tracker.ra_coord[3] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$98.C[3] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$98.C[3] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR(\uut.vga_h_pixel_tracker.o_reset_counter ),
    .O(\uut.vga_h_pixel_tracker.ra_coord[3] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$98.C[4] )
  );
  (* src="top.v:60|../../../lib/interface/Vga.v:88|../../../lib/interface/Vga.v:42|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:60|../../../lib/interface/Vga.v:88|../../../lib/interface/Vga.v:44|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst45 (
    .I0($false),
    .I1($false),
    .I2(\uut.vga_h_pixel_tracker.ra_coord[4] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$98.C[4] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$98.C[4] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR(\uut.vga_h_pixel_tracker.o_reset_counter ),
    .O(\uut.vga_h_pixel_tracker.ra_coord[4] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$98.C[5] )
  );
  (* src="top.v:60|../../../lib/interface/Vga.v:88|../../../lib/interface/Vga.v:42|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:60|../../../lib/interface/Vga.v:88|../../../lib/interface/Vga.v:44|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst46 (
    .I0($false),
    .I1($false),
    .I2(\uut.vga_h_pixel_tracker.ra_coord[5] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$98.C[5] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$98.C[5] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR(\uut.vga_h_pixel_tracker.o_reset_counter ),
    .O(\uut.vga_h_pixel_tracker.ra_coord[5] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$98.C[6] )
  );
  (* src="top.v:60|../../../lib/interface/Vga.v:88|../../../lib/interface/Vga.v:42|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:60|../../../lib/interface/Vga.v:88|../../../lib/interface/Vga.v:44|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst47 (
    .I0($false),
    .I1($false),
    .I2(\uut.vga_h_pixel_tracker.ra_coord[6] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$98.C[6] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$98.C[6] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR(\uut.vga_h_pixel_tracker.o_reset_counter ),
    .O(\uut.vga_h_pixel_tracker.ra_coord[6] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$98.C[7] )
  );
  (* src="top.v:60|../../../lib/interface/Vga.v:88|../../../lib/interface/Vga.v:42|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:60|../../../lib/interface/Vga.v:88|../../../lib/interface/Vga.v:44|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst48 (
    .I0($false),
    .I1($false),
    .I2(\uut.vga_h_pixel_tracker.ra_coord[7] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$98.C[7] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$98.C[7] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR(\uut.vga_h_pixel_tracker.o_reset_counter ),
    .O(\uut.vga_h_pixel_tracker.ra_coord[7] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$98.C[8] )
  );
  (* src="top.v:60|../../../lib/interface/Vga.v:88|../../../lib/interface/Vga.v:42|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:60|../../../lib/interface/Vga.v:88|../../../lib/interface/Vga.v:44|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst49 (
    .I0($false),
    .I1($false),
    .I2(\uut.vga_h_pixel_tracker.ra_coord[8] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$98.C[8] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$98.C[8] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR(\uut.vga_h_pixel_tracker.o_reset_counter ),
    .O(\uut.vga_h_pixel_tracker.ra_coord[8] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$98.C[9] )
  );
  (* src="top.v:60|../../../lib/interface/Vga.v:88|../../../lib/interface/Vga.v:42|/usr/bin/../share/yosys/ice40/cells_map.v:2|top.v:60|../../../lib/interface/Vga.v:88|../../../lib/interface/Vga.v:44|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst50 (
    .I0($false),
    .I1($false),
    .I2(\uut.vga_h_pixel_tracker.ra_coord[9] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$98.C[9] ),
    .CLK(CLK$2),
    .CEN($true),
    .SR(\uut.vga_h_pixel_tracker.o_reset_counter ),
    .O(\uut.vga_h_pixel_tracker.ra_coord[9] )
  );
  (* src="top.v:60|../../../lib/interface/Vga.v:88|../../../lib/interface/Vga.v:42|/usr/bin/../share/yosys/ice40/cells_map.v:2|/usr/bin/../share/yosys/ice40/cells_map.v:44" *)
  ICESTORM_LC #(
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(4'b1001)
  ) $inst51 (
    .I0($abc$1026$new_n103_),
    .I1(\uut.vga_h_pixel_tracker.ra_state[0] ),
    .I2($false),
    .I3($false),
    .CLK(CLK$2),
    .CEN($true),
    .SR($false),
    .O(\uut.vga_h_pixel_tracker.ra_state[0] )
  );
  (* src="top.v:60|../../../lib/interface/Vga.v:88|../../../lib/interface/Vga.v:42|/usr/bin/../share/yosys/ice40/cells_map.v:2|/usr/bin/../share/yosys/ice40/cells_map.v:48" *)
  ICESTORM_LC #(
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(8'b10110100)
  ) $inst52 (
    .I0($abc$1026$new_n103_),
    .I1(\uut.vga_h_pixel_tracker.ra_state[0] ),
    .I2(\uut.vga_h_pixel_tracker.ra_state[1] ),
    .I3($false),
    .CLK(CLK$2),
    .CEN($true),
    .SR($false),
    .O(\uut.vga_h_pixel_tracker.ra_state[1] )
  );
  (* src="top.v:60|../../../lib/interface/Vga.v:107|../../../lib/interface/Vga.v:42|/usr/bin/../share/yosys/ice40/cells_map.v:8|/usr/bin/../share/yosys/ice40/cells_map.v:48" *)
  ICESTORM_LC #(
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(8'b01001011)
  ) $inst53 (
    .I0($abc$1026$new_n98_),
    .I1($abc$1026$new_n97_),
    .I2(\uut.vga_v_pixel_tracker.ra_state[0] ),
    .I3($false),
    .CLK(CLK$2),
    .CEN(\uut.vga_h_pixel_tracker.o_reset_counter ),
    .SR($false),
    .O(\uut.vga_v_pixel_tracker.ra_state[0] )
  );
  (* src="top.v:60|../../../lib/interface/Vga.v:107|../../../lib/interface/Vga.v:42|/usr/bin/../share/yosys/ice40/cells_map.v:8|/usr/bin/../share/yosys/ice40/cells_map.v:52" *)
  ICESTORM_LC #(
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0010111111010000)
  ) $inst54 (
    .I0($abc$1026$new_n97_),
    .I1($abc$1026$new_n98_),
    .I2(\uut.vga_v_pixel_tracker.ra_state[0] ),
    .I3(\uut.vga_v_pixel_tracker.ra_state[1] ),
    .CLK(CLK$2),
    .CEN(\uut.vga_h_pixel_tracker.o_reset_counter ),
    .SR($false),
    .O(\uut.vga_v_pixel_tracker.ra_state[1] )
  );
  (* src="top.v:60|../../../lib/interface/Vga.v:107|../../../lib/interface/Vga.v:42|/usr/bin/../share/yosys/ice40/cells_map.v:8|top.v:60|../../../lib/interface/Vga.v:107|../../../lib/interface/Vga.v:44|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0101101010100101)
  ) $inst55 (
    .I0($false),
    .I1($false),
    .I2(\uut.vga_v_pixel_tracker.ra_coord[0] ),
    .I3($false),
    .CLK(CLK$2),
    .CEN(\uut.vga_h_pixel_tracker.o_reset_counter ),
    .SR(\uut.vga_v_pixel_tracker.o_reset_counter ),
    .O(\uut.vga_v_pixel_tracker.ra_coord[0] )
  );
  (* src="top.v:60|../../../lib/interface/Vga.v:107|../../../lib/interface/Vga.v:42|/usr/bin/../share/yosys/ice40/cells_map.v:8|/usr/bin/../share/yosys/ice40/cells_map.v:40" *)
  ICESTORM_LC #(
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(2'b01)
  ) $inst56 (
    .I0(\uut.vga_v_pixel_tracker.ra_coord[1] ),
    .I1($false),
    .I2($false),
    .I3($false),
    .CLK(CLK$2),
    .CEN(\$abc$1026$auto$dff2dffe.cc:175:make_patterns_logic$868 ),
    .SR(\uut.vga_v_pixel_tracker.o_reset_counter ),
    .O(\uut.vga_v_pixel_tracker.ra_coord[1] )
  );
  (* src="top.v:60|../../../lib/interface/Vga.v:107|../../../lib/interface/Vga.v:42|/usr/bin/../share/yosys/ice40/cells_map.v:8|top.v:60|../../../lib/interface/Vga.v:107|../../../lib/interface/Vga.v:44|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst57 (
    .I0($false),
    .I1($false),
    .I2(\uut.vga_v_pixel_tracker.ra_coord[2] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$104.C[2] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$104.C[2] ),
    .CLK(CLK$2),
    .CEN(\uut.vga_h_pixel_tracker.o_reset_counter ),
    .SR(\uut.vga_v_pixel_tracker.o_reset_counter ),
    .O(\uut.vga_v_pixel_tracker.ra_coord[2] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$104.C[3] )
  );
  (* src="top.v:60|../../../lib/interface/Vga.v:107|../../../lib/interface/Vga.v:42|/usr/bin/../share/yosys/ice40/cells_map.v:8|top.v:60|../../../lib/interface/Vga.v:107|../../../lib/interface/Vga.v:44|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst58 (
    .I0($false),
    .I1($false),
    .I2(\uut.vga_v_pixel_tracker.ra_coord[3] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$104.C[3] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$104.C[3] ),
    .CLK(CLK$2),
    .CEN(\uut.vga_h_pixel_tracker.o_reset_counter ),
    .SR(\uut.vga_v_pixel_tracker.o_reset_counter ),
    .O(\uut.vga_v_pixel_tracker.ra_coord[3] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$104.C[4] )
  );
  (* src="top.v:60|../../../lib/interface/Vga.v:107|../../../lib/interface/Vga.v:42|/usr/bin/../share/yosys/ice40/cells_map.v:8|top.v:60|../../../lib/interface/Vga.v:107|../../../lib/interface/Vga.v:44|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst59 (
    .I0($false),
    .I1($false),
    .I2(\uut.vga_v_pixel_tracker.ra_coord[4] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$104.C[4] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$104.C[4] ),
    .CLK(CLK$2),
    .CEN(\uut.vga_h_pixel_tracker.o_reset_counter ),
    .SR(\uut.vga_v_pixel_tracker.o_reset_counter ),
    .O(\uut.vga_v_pixel_tracker.ra_coord[4] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$104.C[5] )
  );
  (* src="top.v:60|../../../lib/interface/Vga.v:107|../../../lib/interface/Vga.v:42|/usr/bin/../share/yosys/ice40/cells_map.v:8|top.v:60|../../../lib/interface/Vga.v:107|../../../lib/interface/Vga.v:44|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst60 (
    .I0($false),
    .I1($false),
    .I2(\uut.vga_v_pixel_tracker.ra_coord[5] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$104.C[5] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$104.C[5] ),
    .CLK(CLK$2),
    .CEN(\uut.vga_h_pixel_tracker.o_reset_counter ),
    .SR(\uut.vga_v_pixel_tracker.o_reset_counter ),
    .O(\uut.vga_v_pixel_tracker.ra_coord[5] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$104.C[6] )
  );
  (* src="top.v:60|../../../lib/interface/Vga.v:107|../../../lib/interface/Vga.v:42|/usr/bin/../share/yosys/ice40/cells_map.v:8|top.v:60|../../../lib/interface/Vga.v:107|../../../lib/interface/Vga.v:44|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst61 (
    .I0($false),
    .I1($false),
    .I2(\uut.vga_v_pixel_tracker.ra_coord[6] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$104.C[6] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$104.C[6] ),
    .CLK(CLK$2),
    .CEN(\uut.vga_h_pixel_tracker.o_reset_counter ),
    .SR(\uut.vga_v_pixel_tracker.o_reset_counter ),
    .O(\uut.vga_v_pixel_tracker.ra_coord[6] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$104.C[7] )
  );
  (* src="top.v:60|../../../lib/interface/Vga.v:107|../../../lib/interface/Vga.v:42|/usr/bin/../share/yosys/ice40/cells_map.v:8|top.v:60|../../../lib/interface/Vga.v:107|../../../lib/interface/Vga.v:44|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst62 (
    .I0($false),
    .I1($false),
    .I2(\uut.vga_v_pixel_tracker.ra_coord[7] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$104.C[7] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$104.C[7] ),
    .CLK(CLK$2),
    .CEN(\uut.vga_h_pixel_tracker.o_reset_counter ),
    .SR(\uut.vga_v_pixel_tracker.o_reset_counter ),
    .O(\uut.vga_v_pixel_tracker.ra_coord[7] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$104.C[8] )
  );
  (* src="top.v:60|../../../lib/interface/Vga.v:107|../../../lib/interface/Vga.v:42|/usr/bin/../share/yosys/ice40/cells_map.v:8|top.v:60|../../../lib/interface/Vga.v:107|../../../lib/interface/Vga.v:44|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst63 (
    .I0($false),
    .I1($false),
    .I2(\uut.vga_v_pixel_tracker.ra_coord[8] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$104.C[8] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$104.C[8] ),
    .CLK(CLK$2),
    .CEN(\uut.vga_h_pixel_tracker.o_reset_counter ),
    .SR(\uut.vga_v_pixel_tracker.o_reset_counter ),
    .O(\uut.vga_v_pixel_tracker.ra_coord[8] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$104.C[9] )
  );
  (* src="top.v:60|../../../lib/interface/Vga.v:107|../../../lib/interface/Vga.v:42|/usr/bin/../share/yosys/ice40/cells_map.v:8|top.v:60|../../../lib/interface/Vga.v:107|../../../lib/interface/Vga.v:44|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .DFF_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst64 (
    .I0($false),
    .I1($false),
    .I2(\uut.vga_v_pixel_tracker.ra_coord[9] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$104.C[9] ),
    .CLK(CLK$2),
    .CEN(\uut.vga_h_pixel_tracker.o_reset_counter ),
    .SR(\uut.vga_v_pixel_tracker.o_reset_counter ),
    .O(\uut.vga_v_pixel_tracker.ra_coord[9] )
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:52" *)
  ICESTORM_LC #(
    .LUT_INIT(16'b0100000000000000)
  ) $inst65 (
    .I0(\uut.vga_h_pixel_tracker.ra_coord[5] ),
    .I1(\$abc$1026$auto$simplemap.cc:127:simplemap_reduce$263[0]_new_inv_ ),
    .I2($abc$1026$new_n69_),
    .I3(\uut.vga_h_pixel_tracker.ra_coord[4] ),
    .O(\uut.vga_h_pixel_tracker.o_reset_counter )
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:52" *)
  ICESTORM_LC #(
    .LUT_INIT(16'b0001000000000000)
  ) $inst66 (
    .I0(\uut.vga_h_pixel_tracker.ra_coord[6] ),
    .I1(\uut.vga_h_pixel_tracker.ra_coord[7] ),
    .I2(\uut.vga_h_pixel_tracker.ra_coord[8] ),
    .I3(\uut.vga_h_pixel_tracker.ra_coord[9] ),
    .O($abc$1026$new_n69_)
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:52" *)
  ICESTORM_LC #(
    .LUT_INIT(16'b1000000000000000)
  ) $inst67 (
    .I0(\uut.vga_h_pixel_tracker.ra_coord[1] ),
    .I1(\uut.vga_h_pixel_tracker.ra_coord[2] ),
    .I2(\uut.vga_h_pixel_tracker.ra_coord[3] ),
    .I3(\uut.vga_h_pixel_tracker.ra_coord[0] ),
    .O(\$abc$1026$auto$simplemap.cc:127:simplemap_reduce$263[0]_new_inv_ )
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:52" *)
  ICESTORM_LC #(
    .LUT_INIT(16'b0100000000000000)
  ) $inst68 (
    .I0(\uut.vga_v_pixel_tracker.ra_coord[1] ),
    .I1($abc$1026$new_n72_),
    .I2(\uut.vga_v_pixel_tracker.ra_coord[2] ),
    .I3(\uut.vga_v_pixel_tracker.ra_coord[3] ),
    .O(\uut.vga_v_pixel_tracker.o_reset_counter )
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:52" *)
  ICESTORM_LC #(
    .LUT_INIT(16'b0001000000000000)
  ) $inst69 (
    .I0(\uut.vga_v_pixel_tracker.ra_coord[6] ),
    .I1(\uut.vga_v_pixel_tracker.ra_coord[7] ),
    .I2($abc$1026$new_n73_),
    .I3(\uut.vga_v_pixel_tracker.ra_coord[9] ),
    .O($abc$1026$new_n72_)
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:52" *)
  ICESTORM_LC #(
    .LUT_INIT(16'b0000000000000001)
  ) $inst70 (
    .I0(\uut.vga_v_pixel_tracker.ra_coord[0] ),
    .I1(\uut.vga_v_pixel_tracker.ra_coord[8] ),
    .I2(\uut.vga_v_pixel_tracker.ra_coord[4] ),
    .I3(\uut.vga_v_pixel_tracker.ra_coord[5] ),
    .O($abc$1026$new_n73_)
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:48" *)
  ICESTORM_LC #(
    .LUT_INIT(8'b11100000)
  ) $inst71 (
    .I0(\uut.vga_v_pixel_tracker.ra_coord[0] ),
    .I1(\uut.vga_v_pixel_tracker.o_reset_counter ),
    .I2(\uut.vga_h_pixel_tracker.o_reset_counter ),
    .I3($false),
    .O(\$abc$1026$auto$dff2dffe.cc:175:make_patterns_logic$868 )
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:44" *)
  ICESTORM_LC #(
    .LUT_INIT(4'b1000)
  ) $inst72 (
    .I0($abc$1026$visible_new_),
    .I1(\in_r[0] ),
    .I2($false),
    .I3($false),
    .O(VGA_R0$2)
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:52" *)
  ICESTORM_LC #(
    .LUT_INIT(16'b0000000000000001)
  ) $inst73 (
    .I0(\uut.vga_h_pixel_tracker.ra_state[0] ),
    .I1(\uut.vga_h_pixel_tracker.ra_state[1] ),
    .I2(\uut.vga_v_pixel_tracker.ra_state[0] ),
    .I3(\uut.vga_v_pixel_tracker.ra_state[1] ),
    .O($abc$1026$visible_new_)
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:44" *)
  ICESTORM_LC #(
    .LUT_INIT(4'b1000)
  ) $inst74 (
    .I0($abc$1026$visible_new_),
    .I1(\in_r[1] ),
    .I2($false),
    .I3($false),
    .O(VGA_R1$2)
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:44" *)
  ICESTORM_LC #(
    .LUT_INIT(4'b1000)
  ) $inst75 (
    .I0($abc$1026$visible_new_),
    .I1(\in_r[2] ),
    .I2($false),
    .I3($false),
    .O(VGA_R2$2)
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:44" *)
  ICESTORM_LC #(
    .LUT_INIT(4'b1000)
  ) $inst76 (
    .I0($abc$1026$visible_new_),
    .I1(\in_g[0] ),
    .I2($false),
    .I3($false),
    .O(VGA_G0$2)
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:44" *)
  ICESTORM_LC #(
    .LUT_INIT(4'b1000)
  ) $inst77 (
    .I0($abc$1026$visible_new_),
    .I1(\in_g[1] ),
    .I2($false),
    .I3($false),
    .O(VGA_G1$2)
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:44" *)
  ICESTORM_LC #(
    .LUT_INIT(4'b1000)
  ) $inst78 (
    .I0($abc$1026$visible_new_),
    .I1(\in_g[2] ),
    .I2($false),
    .I3($false),
    .O(VGA_G2$2)
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:44" *)
  ICESTORM_LC #(
    .LUT_INIT(4'b1000)
  ) $inst79 (
    .I0($abc$1026$visible_new_),
    .I1(\in_b[0] ),
    .I2($false),
    .I3($false),
    .O(VGA_B0$2)
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:44" *)
  ICESTORM_LC #(
    .LUT_INIT(4'b1000)
  ) $inst80 (
    .I0($abc$1026$visible_new_),
    .I1(\in_b[1] ),
    .I2($false),
    .I3($false),
    .O(VGA_B1$2)
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:44" *)
  ICESTORM_LC #(
    .LUT_INIT(4'b1000)
  ) $inst81 (
    .I0($abc$1026$visible_new_),
    .I1(\in_b[2] ),
    .I2($false),
    .I3($false),
    .O(VGA_B2$2)
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:44" *)
  ICESTORM_LC #(
    .LUT_INIT(4'b0100)
  ) $inst82 (
    .I0(\uut.vga_v_pixel_tracker.ra_state[0] ),
    .I1(\uut.vga_v_pixel_tracker.ra_state[1] ),
    .I2($false),
    .I3($false),
    .O(VGA_VS$2)
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:44" *)
  ICESTORM_LC #(
    .LUT_INIT(4'b0100)
  ) $inst83 (
    .I0(\uut.vga_h_pixel_tracker.ra_state[0] ),
    .I1(\uut.vga_h_pixel_tracker.ra_state[1] ),
    .I2($false),
    .I3($false),
    .O(VGA_HS$2)
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:44" *)
  ICESTORM_LC #(
    .LUT_INIT(4'b0110)
  ) $inst84 (
    .I0(\uut.vga_v_pixel_tracker.ra_coord[0] ),
    .I1(\uut.vga_h_pixel_tracker.ra_coord[0] ),
    .I2($false),
    .I3($false),
    .O(\$abc$1026$auto$alumacc.cc:474:replace_alu$92.BB[0] )
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:44" *)
  ICESTORM_LC #(
    .LUT_INIT(4'b0110)
  ) $inst85 (
    .I0(\uut.vga_h_pixel_tracker.ra_coord[1] ),
    .I1(\uut.vga_v_pixel_tracker.ra_coord[1] ),
    .I2($false),
    .I3($false),
    .O(\$abc$1026$auto$alumacc.cc:474:replace_alu$92.BB[1] )
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:44" *)
  ICESTORM_LC #(
    .LUT_INIT(4'b0110)
  ) $inst86 (
    .I0(\uut.vga_h_pixel_tracker.ra_coord[2] ),
    .I1(\uut.vga_v_pixel_tracker.ra_coord[2] ),
    .I2($false),
    .I3($false),
    .O(\$abc$1026$auto$alumacc.cc:474:replace_alu$92.BB[2] )
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:44" *)
  ICESTORM_LC #(
    .LUT_INIT(4'b0110)
  ) $inst87 (
    .I0(\uut.vga_h_pixel_tracker.ra_coord[3] ),
    .I1(\uut.vga_v_pixel_tracker.ra_coord[3] ),
    .I2($false),
    .I3($false),
    .O(\$abc$1026$auto$alumacc.cc:474:replace_alu$92.BB[3] )
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:44" *)
  ICESTORM_LC #(
    .LUT_INIT(4'b0110)
  ) $inst88 (
    .I0(\uut.vga_h_pixel_tracker.ra_coord[4] ),
    .I1(\uut.vga_v_pixel_tracker.ra_coord[4] ),
    .I2($false),
    .I3($false),
    .O(\$abc$1026$auto$alumacc.cc:474:replace_alu$92.BB[4] )
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:44" *)
  ICESTORM_LC #(
    .LUT_INIT(4'b0110)
  ) $inst89 (
    .I0(\uut.vga_h_pixel_tracker.ra_coord[5] ),
    .I1(\uut.vga_v_pixel_tracker.ra_coord[5] ),
    .I2($false),
    .I3($false),
    .O(\$abc$1026$auto$alumacc.cc:474:replace_alu$92.BB[5] )
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:44" *)
  ICESTORM_LC #(
    .LUT_INIT(4'b0110)
  ) $inst90 (
    .I0(\uut.vga_h_pixel_tracker.ra_coord[6] ),
    .I1(\uut.vga_v_pixel_tracker.ra_coord[6] ),
    .I2($false),
    .I3($false),
    .O(\$abc$1026$auto$alumacc.cc:474:replace_alu$92.BB[6] )
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:44" *)
  ICESTORM_LC #(
    .LUT_INIT(4'b0110)
  ) $inst91 (
    .I0(\uut.vga_h_pixel_tracker.ra_coord[7] ),
    .I1(\uut.vga_v_pixel_tracker.ra_coord[7] ),
    .I2($false),
    .I3($false),
    .O(\$abc$1026$auto$alumacc.cc:474:replace_alu$92.BB[7] )
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:44" *)
  ICESTORM_LC #(
    .LUT_INIT(4'b0110)
  ) $inst92 (
    .I0(\uut.vga_h_pixel_tracker.ra_coord[8] ),
    .I1(\uut.vga_v_pixel_tracker.ra_coord[8] ),
    .I2($false),
    .I3($false),
    .O(\$abc$1026$auto$alumacc.cc:474:replace_alu$92.BB[8] )
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:52" *)
  ICESTORM_LC #(
    .LUT_INIT(16'b1011110011111111)
  ) $inst93 (
    .I0(\uut.vga_v_pixel_tracker.ra_coord[1] ),
    .I1(\uut.vga_v_pixel_tracker.ra_coord[2] ),
    .I2(\uut.vga_v_pixel_tracker.ra_coord[3] ),
    .I3($abc$1026$new_n72_),
    .O($abc$1026$new_n97_)
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:52" *)
  ICESTORM_LC #(
    .LUT_INIT(16'b1000000000000000)
  ) $inst94 (
    .I0($abc$1026$new_n99_),
    .I1($abc$1026$new_n100_),
    .I2(\uut.vga_v_pixel_tracker.ra_coord[2] ),
    .I3(\uut.vga_v_pixel_tracker.ra_coord[3] ),
    .O($abc$1026$new_n98_)
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:52" *)
  ICESTORM_LC #(
    .LUT_INIT(16'b0001000000000000)
  ) $inst95 (
    .I0(\uut.vga_v_pixel_tracker.ra_coord[5] ),
    .I1(\uut.vga_v_pixel_tracker.ra_coord[9] ),
    .I2(\uut.vga_v_pixel_tracker.ra_coord[7] ),
    .I3(\uut.vga_v_pixel_tracker.ra_coord[6] ),
    .O($abc$1026$new_n99_)
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:52" *)
  ICESTORM_LC #(
    .LUT_INIT(16'b1000000000000000)
  ) $inst96 (
    .I0(\uut.vga_v_pixel_tracker.ra_coord[0] ),
    .I1(\uut.vga_v_pixel_tracker.ra_coord[8] ),
    .I2(\uut.vga_v_pixel_tracker.ra_coord[1] ),
    .I3(\uut.vga_v_pixel_tracker.ra_coord[4] ),
    .O($abc$1026$new_n100_)
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:52" *)
  ICESTORM_LC #(
    .LUT_INIT(16'b0000000000001101)
  ) $inst97 (
    .I0($abc$1026$new_n110_),
    .I1($abc$1026$new_n118_),
    .I2($abc$1026$new_n108_),
    .I3(\uut.vga_h_pixel_tracker.o_reset_counter ),
    .O($abc$1026$new_n103_)
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:44" *)
  ICESTORM_LC #(
    .LUT_INIT(4'b0100)
  ) $inst98 (
    .I0(\uut.vga_h_pixel_tracker.ra_coord[1] ),
    .I1(\uut.vga_h_pixel_tracker.ra_coord[0] ),
    .I2($false),
    .I3($false),
    .O(\$abc$1026$auto$simplemap.cc:127:simplemap_reduce$310[0]_new_inv_ )
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:48" *)
  ICESTORM_LC #(
    .LUT_INIT(8'b10000000)
  ) $inst99 (
    .I0($abc$1026$new_n69_),
    .I1(\$abc$1026$auto$simplemap.cc:127:simplemap_reduce$310[0]_new_inv_ ),
    .I2($abc$1026$new_n109_),
    .I3($false),
    .O($abc$1026$new_n108_)
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:52" *)
  ICESTORM_LC #(
    .LUT_INIT(16'b0001000000000000)
  ) $inst100 (
    .I0(\uut.vga_h_pixel_tracker.ra_coord[5] ),
    .I1(\uut.vga_h_pixel_tracker.ra_coord[4] ),
    .I2(\uut.vga_h_pixel_tracker.ra_coord[2] ),
    .I3(\uut.vga_h_pixel_tracker.ra_coord[3] ),
    .O($abc$1026$new_n109_)
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:52" *)
  ICESTORM_LC #(
    .LUT_INIT(16'b0100000000000000)
  ) $inst101 (
    .I0(\uut.vga_h_pixel_tracker.ra_coord[8] ),
    .I1(\uut.vga_h_pixel_tracker.ra_coord[4] ),
    .I2(\uut.vga_h_pixel_tracker.ra_coord[5] ),
    .I3(\uut.vga_h_pixel_tracker.ra_coord[9] ),
    .O($abc$1026$new_n110_)
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:52" *)
  ICESTORM_LC #(
    .LUT_INIT(16'b0000000111110000)
  ) $inst102 (
    .I0(\uut.vga_h_pixel_tracker.ra_coord[2] ),
    .I1(\uut.vga_h_pixel_tracker.ra_coord[3] ),
    .I2(\uut.vga_h_pixel_tracker.ra_coord[6] ),
    .I3(\uut.vga_h_pixel_tracker.ra_coord[7] ),
    .O($abc$1026$new_n117_)
  );
  (* src="/usr/bin/../share/yosys/ice40/cells_map.v:52" *)
  ICESTORM_LC #(
    .LUT_INIT(16'b0011010111111111)
  ) $inst103 (
    .I0(\$abc$1026$auto$simplemap.cc:127:simplemap_reduce$310[0]_new_inv_ ),
    .I1(\$abc$1026$auto$simplemap.cc:127:simplemap_reduce$263[0]_new_inv_ ),
    .I2(\uut.vga_h_pixel_tracker.ra_coord[6] ),
    .I3($abc$1026$new_n117_),
    .O($abc$1026$new_n118_)
  );
  (* src="top.v:54|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .LUT_INIT(16'b0110100110010110)
  ) $inst104 (
    .I0($false),
    .I1(\ra_time[20] ),
    .I2(\$abc$1026$auto$alumacc.cc:474:replace_alu$92.BB[0] ),
    .I3($false),
    .O(\in_b[0] )
  );
  (* src="top.v:54|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst105 (
    .I0($false),
    .I1(\ra_time[21] ),
    .I2(\$abc$1026$auto$alumacc.cc:474:replace_alu$92.BB[1] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$92.C[1] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$92.C[1] ),
    .O(\in_b[1] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$92.C[2] )
  );
  (* src="top.v:54|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst106 (
    .I0($false),
    .I1(\ra_time[22] ),
    .I2(\$abc$1026$auto$alumacc.cc:474:replace_alu$92.BB[2] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$92.C[2] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$92.C[2] ),
    .O(\in_b[2] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$92.C[3] )
  );
  (* src="top.v:54|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst107 (
    .I0($false),
    .I1(\ra_time[23] ),
    .I2(\$abc$1026$auto$alumacc.cc:474:replace_alu$92.BB[3] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$92.C[3] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$92.C[3] ),
    .O(\in_g[0] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$92.C[4] )
  );
  (* src="top.v:54|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst108 (
    .I0($false),
    .I1(\ra_time[24] ),
    .I2(\$abc$1026$auto$alumacc.cc:474:replace_alu$92.BB[4] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$92.C[4] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$92.C[4] ),
    .O(\in_g[1] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$92.C[5] )
  );
  (* src="top.v:54|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst109 (
    .I0($false),
    .I1(\ra_time[25] ),
    .I2(\$abc$1026$auto$alumacc.cc:474:replace_alu$92.BB[5] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$92.C[5] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$92.C[5] ),
    .O(\in_g[2] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$92.C[6] )
  );
  (* src="top.v:54|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst110 (
    .I0($false),
    .I1(\ra_time[26] ),
    .I2(\$abc$1026$auto$alumacc.cc:474:replace_alu$92.BB[6] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$92.C[6] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$92.C[6] ),
    .O(\in_r[0] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$92.C[7] )
  );
  (* src="top.v:54|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1), 
    .LUT_INIT(16'b0110100110010110)
  ) $inst111 (
    .I0($false),
    .I1(\ra_time[27] ),
    .I2(\$abc$1026$auto$alumacc.cc:474:replace_alu$92.BB[7] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$92.C[7] ),
    .CIN(\$auto$alumacc.cc:474:replace_alu$92.C[7] ),
    .O(\in_r[1] ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$92.C[8] )
  );
  (* src="top.v:54|/usr/bin/../share/yosys/ice40/arith_map.v:53" *)
  ICESTORM_LC #(
    .LUT_INIT(16'b0110100110010110)
  ) $inst112 (
    .I0($false),
    .I1(\ra_time[28] ),
    .I2(\$abc$1026$auto$alumacc.cc:474:replace_alu$92.BB[8] ),
    .I3(\$auto$alumacc.cc:474:replace_alu$92.C[8] ),
    .O(\in_r[2] )
  );
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1)
  ) $inst113 (
    .I0($false),
    .I1(\uut.vga_v_pixel_tracker.ra_coord[0] ),
    .I2($false),
    .I3($false),
    .CIN($true),
    .COUT(\uut.vga_v_pixel_tracker.ra_coord[0]$2 )
  );
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1)
  ) $inst114 (
    .I1($false),
    .I2(\uut.vga_v_pixel_tracker.ra_coord[1] ),
    .CIN(\uut.vga_v_pixel_tracker.ra_coord[0]$2 ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$104.C[2] )
  );
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1)
  ) $inst115 (
    .I1(\ra_time[20] ),
    .I2(\$abc$1026$auto$alumacc.cc:474:replace_alu$92.BB[0] ),
    .CIN($false),
    .COUT(\$auto$alumacc.cc:474:replace_alu$92.C[1] )
  );
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1)
  ) $inst116 (
    .I0($false),
    .I1(\ra_time[0] ),
    .I2($false),
    .I3($false),
    .CIN($true),
    .COUT(\ra_time[0]$2 )
  );
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1)
  ) $inst117 (
    .I1($false),
    .I2(\ra_time[1] ),
    .CIN(\ra_time[0]$2 ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$95.C[2] )
  );
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1)
  ) $inst118 (
    .I0($false),
    .I1(\uut.vga_h_pixel_tracker.ra_coord[0] ),
    .I2($false),
    .I3($false),
    .CIN($true),
    .COUT(\uut.vga_h_pixel_tracker.ra_coord[0]$2 )
  );
  ICESTORM_LC #(
    .CARRY_ENABLE(1'b1)
  ) $inst119 (
    .I1($false),
    .I2(\uut.vga_h_pixel_tracker.ra_coord[1] ),
    .CIN(\uut.vga_h_pixel_tracker.ra_coord[0]$2 ),
    .COUT(\$auto$alumacc.cc:474:replace_alu$98.C[2] )
  );
endmodule
