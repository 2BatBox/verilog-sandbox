module SyncChain_tb();
endmodule
