module Dummy();
endmodule
